CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 100 10
176 80 1278 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
11
2 +V
167 150 156 0 1 3
0 4
0
0 0 54240 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 1025 133 0 17 19
10 11 10 9 8 7 6 5 18 2
1 1 0 1 1 0 1 2
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
391 0 0
2
5.89883e-315 0
0
7 Ground~
168 982 78 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3124 0 0
2
5.89883e-315 0
0
7 Pulser~
4 131 390 0 10 12
0 19 20 3 3 0 0 5 5 1
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3421 0 0
2
5.89883e-315 0
0
6 74112~
219 383 269 0 7 32
0 4 17 3 17 4 21 16
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 4 0
1 U
8157 0 0
2
5.89883e-315 0
0
6 74LS48
188 862 370 0 14 29
0 12 14 16 17 22 23 5 6 7
8 9 10 11 24
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
5572 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 694 106 0 3 22
0 15 14 13
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 487 105 0 3 22
0 17 16 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
5.89883e-315 0
0
6 74112~
219 775 263 0 7 32
0 4 13 3 13 4 25 12
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
4747 0 0
2
5.89883e-315 0
0
6 74112~
219 569 267 0 7 32
0 4 15 3 15 4 26 14
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
972 0 0
2
5.89883e-315 0
0
6 74112~
219 197 269 0 7 32
0 4 4 3 4 4 27 17
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3472 0 0
2
5.89883e-315 0
0
38
4 0 3 0 0 4096 0 4 0 0 2 3
161 390
161 381
159 381
3 0 3 0 0 8192 0 4 0 0 35 3
155 381
169 381
169 323
5 0 4 0 0 4096 0 10 0 0 10 2
569 279
569 297
5 0 4 0 0 0 0 5 0 0 10 2
383 281
383 297
1 0 4 0 0 0 0 5 0 0 9 2
383 206
383 192
1 0 4 0 0 0 0 10 0 0 9 2
569 204
569 192
1 0 4 0 0 0 0 11 0 0 9 2
197 206
197 192
0 0 4 0 0 4096 0 0 0 9 10 2
287 192
287 297
0 1 4 0 0 4224 0 0 9 11 0 3
150 192
775 192
775 200
5 5 4 0 0 0 0 11 9 0 0 4
197 281
197 297
775 297
775 275
1 0 4 0 0 0 0 1 0 0 12 2
150 165
150 233
0 2 4 0 0 0 0 0 11 13 0 2
150 233
173 233
4 2 4 0 0 0 0 11 11 0 0 4
173 251
149 251
149 233
173 233
9 1 2 0 0 4112 0 2 3 0 0 4
1025 91
1025 68
982 68
982 72
7 7 5 0 0 8320 0 6 2 0 0 3
894 334
1040 334
1040 169
8 6 6 0 0 8320 0 6 2 0 0 3
894 343
1034 343
1034 169
9 5 7 0 0 8320 0 6 2 0 0 3
894 352
1028 352
1028 169
10 4 8 0 0 8320 0 6 2 0 0 3
894 361
1022 361
1022 169
11 3 9 0 0 8320 0 6 2 0 0 3
894 370
1016 370
1016 169
12 2 10 0 0 8320 0 6 2 0 0 3
894 379
1010 379
1010 169
13 1 11 0 0 8320 0 6 2 0 0 3
894 388
1004 388
1004 169
7 1 12 0 0 8320 0 9 6 0 0 4
799 227
811 227
811 334
830 334
4 0 13 0 0 4096 0 9 0 0 24 3
751 245
720 245
720 227
2 3 13 0 0 8320 0 9 7 0 0 4
751 227
719 227
719 106
715 106
0 2 14 0 0 8320 0 0 6 26 0 3
657 231
657 343
830 343
7 2 14 0 0 0 0 10 7 0 0 4
593 231
658 231
658 115
670 115
4 0 15 0 0 8192 0 10 0 0 28 3
545 249
536 249
536 231
2 0 15 0 0 8192 0 10 0 0 29 3
545 231
522 231
522 105
3 1 15 0 0 8320 0 8 7 0 0 4
508 105
522 105
522 97
670 97
3 0 3 0 0 8192 0 10 0 0 35 3
539 240
529 240
529 323
0 3 16 0 0 8320 0 0 6 32 0 3
461 233
461 352
830 352
7 2 16 0 0 0 0 5 8 0 0 4
407 233
461 233
461 114
463 114
4 0 17 0 0 4096 0 5 0 0 38 3
359 251
319 251
319 233
3 0 3 0 0 0 0 5 0 0 35 3
353 242
349 242
349 323
3 3 3 0 0 12416 0 11 9 0 0 6
167 242
163 242
163 323
737 323
737 236
745 236
0 4 17 0 0 8320 0 0 6 38 0 3
253 233
253 361
830 361
1 0 17 0 0 0 0 8 0 0 33 3
463 96
319 96
319 233
7 2 17 0 0 0 0 11 5 0 0 2
221 233
359 233
2
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
281 33 588 68
291 41 577 64
22 BINARY 4-BIT SYNCHRONO
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
566 33 756 68
576 41 745 64
13 US UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
